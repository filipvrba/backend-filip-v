module server

pub struct Health {
	status_code int
	status string
}
