module cli

import rb

const(
	app_name = rb.get_app_name()
	app_full_name = "Backend-Filip"
	version = '1.0.0'
	path_config = "./shared/config.json"
)