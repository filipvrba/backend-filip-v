module cli

pub struct Cli {
pub:
	arguments Arguments = get_arguments()
}
